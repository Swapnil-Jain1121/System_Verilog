module top ();

  initial begin
    $display("process#1");
  end

  initial begin
    $display("process#2");
  end

  initial begin
    $display("process#3");
  end

  initial begin
    $display("process#4");
  end

endmodule

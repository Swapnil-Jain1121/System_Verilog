class data_pkt extends usb_base_pkt;

  function bit [5:0] calc_crc5();

  endfunction
endclass
